subck 0603C0 0 1 2 3 4

#include NN.subs

TMS:TP0 0 +1 +A1 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT
TMS:TP1 0 +2 -A1 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT

TMS:TP2 0 +4 +B1 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT
TMS:TP3 0 +3 -B1 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT

C:Cp A1 B1 c=0.01e-12

*TMSGAP:TG1 0 A2 B2 M1=TP1 M2=TP2



VIA:V1 0 B1 $DURVIA D=0.5e-3 FOOTPRINT="RPAD=0.01e-3"
C:CC A1 B1 c=100e-12 l=0.75e-9 tand=1e-4 rskin=2.5e-6 ESRF=100e6 ESR=70e-3 $TEMP
func:C1 type=4 v1=39 data=NPO_0603.txt CC:C(1) CC:ESR(2) CC:ESRF(3)

FP:M2PADM:P A1 B1 D=0.9e-3 B=0.6e-3 W=0.9e-3 DIR1=1 DIR2=1 LABEL=C VALUE=CC:C

