subck 0603C0 0 1 2 3
#include NN.subs

TMS:TP0 0 +1  +A1 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT
TMS:TP1 0 +2  -A1 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT

TMS:TP2 0 B1 B2 $DUR len=0.3e-3 w=0.9e-3 FOOTPRINT
TMS:TP3 0 +3 B1 $DUR len=0.3e-3 w=0.9e-3 FOOTPRINT

R:R2 A1 X1 r=1 $TEMP
C:CP X1 XP c=0.1e-12 
R:RP XP B1 r=1 $TEMP
L:LS X1 B1 l=1e-9 rskin=1 $TEMP
 
func:L1 type=4 v1=10 data=IND_0603.txt LS:L(1) RP:R(2) R2:R(3) CP:C(4) LS:RSKIN(5)
**1-48**L, RP, R2, C, rskin@1GHz

FP:M2PADM:P A1 +B1 D=0.9e-3 B=0.6e-3 W=0.9e-3 DIR1=1 DIR2=0 LABEL=L VALUE=LS:L
