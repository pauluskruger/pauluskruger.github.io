subck Sparm S G D

T:TA S G D atf35143b.s2p
.ends