subck ATF35 0 1 2
#include NN.subs


*Gate&Drain pads
TMS:TG1 0 1 G  $DUR len=0.3e-3 w=0.5e-3 FOOTPRINT
TMS:TG2 0 G G1 $DUR len=0.3e-3 w=0.5e-3 FOOTPRINT OPEN=2

TMS:TD1 0 2 D  $DUR len=0.3e-3 w=0.5e-3 FOOTPRINT
TMS:TD2 0 -D D1 $DUR len=0.3e-3 w=0.5e-3 FOOTPRINT OPEN=2

FP:EQ:EQ0 G D X=2.2e-3 Y=0 ANG=0


*Transistor
CKT:T1 sa1 sb1 G D atf35143.ckt
R:RS sa1 0 r=50 $TEMP
*Source footprints
TMS:TSA0 0 -sa sa1 $DUR len=0.45e-3 w=1.0e-3 FOOTPRINT 
TMS:TSA1 0 +sa sa2 $DUR len=0.45e-3 w=1.0e-3 FOOTPRINT
TMS:TSA2 0 sa1 sa0 $DUR len=0.45e-3 w=1.0e-3 FOOTPRINT open=2
TMS:TSA3 0 sa2 sa3 $DUR len=0.45e-3 w=1.0e-3 FOOTPRINT open=2

TMS:TSB0 0 -sb sb1 $DUR len=0.45e-3 w=1.0e-3 FOOTPRINT 
TMS:TSB1 0 +sb sb2 $DUR len=0.45e-3 w=1.0e-3 FOOTPRINT
TMS:TSB2 0 sb1 sb0 $DUR len=0.45e-3 w=1.0e-3 FOOTPRINT open=2
TMS:TSB3 0 sb2 sb3 $DUR len=0.45e-3 w=1.0e-3 FOOTPRINT open=2

FP:EQ:EQ1 G sa1 X=0.6e-3 Y=1.2e-3 ANG=-52
FP:EQ:EQ2 D sb1 X=0.6e-3 Y=1.1e-3 ANG=-52


*Source1 capacitor
C:CS1 sa1 va1 c=100e-12 l=0.75e-9 tand=1e-4 rskin=2.5e-6 ESRF=100e6 ESR=70e-3 $TEMP
func:CS1V type=4 v1=39 data=NPO_0603.txt CS1:C(1) CS1:ESR(2) CS1:ESRF(3)

C:CS2 sa2 va2 c=100e-12 l=0.75e-9 tand=1e-4 rskin=2.5e-6 ESRF=100e6 ESR=70e-3 $TEMP
func:CS2V type=4 v1=39 data=NPO_0603.txt CS2:C(1) CS2:ESR(2) CS2:ESRF(3)

C:CS3 sb1 vb1 c=100e-12 l=0.75e-9 tand=1e-4 rskin=2.5e-6 ESRF=100e6 ESR=70e-3 $TEMP
func:CS3V type=4 v1=39 data=NPO_0603.txt CS3:C(1) CS3:ESR(2) CS3:ESRF(3)

C:CS4 sb2 vb2 c=100e-12 l=0.75e-9 tand=1e-4 rskin=2.5e-6 ESRF=100e6 ESR=70e-3 $TEMP
func:CS4V type=4 v1=39 data=NPO_0603.txt CS4:C(1) CS4:ESR(2) CS4:ESRF(3)
FP:EQ:POFF1 sa saF X=0 Y=-0.2e-3 ANG=0
FP:EQ:POFF2 sb sbF X=0 Y=-0.2e-3 ANG=0
FP:M2PAD:CS1 +saF +va D=0.9e-3 B=0.6e-3 W=0.9e-3 LABEL=C VALUE=CS1:C DIR1=1 DIR2=-1
FP:M2PAD:CS2 -saF -va D=0.9e-3 B=0.6e-3 W=0.9e-3 LABEL=C VALUE=CS2:C DIR1=-1 DIR2=1
FP:M2PAD:CS3 +sbF +vb D=0.9e-3 B=0.6e-3 W=0.9e-3 LABEL=C VALUE=CS1:C DIR1=1 DIR2=-1
FP:M2PAD:CS4 -sbF -vb D=0.9e-3 B=0.6e-3 W=0.9e-3 LABEL=C VALUE=CS2:C DIR1=-1 DIR2=1

TMS:TVA0 0 +va va1 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT 
TMS:TVA1 0 -va va2 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT
TMS:TVA2 0 va1 va0 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT
TMS:TVA3 0 va2 va3 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT

TMS:TVB0 0 +vb vb1 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT 
TMS:TVB1 0 -vb vb2 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT
TMS:TVB2 0 vb1 vb0 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT
TMS:TVB3 0 vb2 vb3 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT

VIA:V1 0 va1 $DURVIA D=0.5e-3 FOOTPRINT="RPAD=0.01e-3"
VIA:V2 0 va2 $DURVIA D=0.5e-3 FOOTPRINT="RPAD=0.01e-3"
VIA:V3 0 vb1 $DURVIA D=0.5e-3 FOOTPRINT="RPAD=0.01e-3"
VIA:V4 0 vb2 $DURVIA D=0.5e-3 FOOTPRINT="RPAD=0.01e-3"

*TMSR:R1 0 sa1 va1 $DURR w=0.9e03 LEN=1.5e-3 R=100
R:RS sa1 va1 r=50 $TEMP

*Drain resistor
*CKT:LD 0 +D 2 0603L0.ckt FOOTPRINT
*CKT:RD 0 +D 2 0603R0.ckt FOOTPRINT
*CKT:RD 0 +D2 D10 0603R0.ckt FOOTPRINT

*TMS:TD3 0 D3 D4  $DUR len=0.5e-3 w=0.2e-3 FOOTPRINT
*TMS:TD4 0 D5 D6  $DUR len=2.1e-3 w=0.2e-3 FOOTPRINT
*TMS:TD5 0 D7 D8  $DUR len=0.5e-3 w=0.2e-3 FOOTPRINT
*TMS:TD6 0 D9 2   $DUR len=0.1e-3 w=0.6e-3 FOOTPRINT

*TMSTEE:TE1 0 +D +D2 +D3 M1=TD2 M2=RD:TP0 M3=TD3 FOOTPRINT
*TMSCNR:TC1 0 D4 D5 $DUR w=0.2e-3 FOOTPRINT
*TMSCNR:TC2 0 D6 D7 $DUR w=0.2e-3 FOOTPRINT
*TMSTEE:TE2 0 -D10 -D9 +D8 M1=RD:TP3 M2=TD6 M3=TD5 FOOTPRINT

*FUNC:FL type=0 v1=0.8e-3 v2=0 TD3:LEN(1,0) TD5:LEN(1,0)
*FUNC:FW type=0 v1=0.3e-3 v2=0 TD3:W(1,0) TD4:W(1,0) TD5:W(1,5) TC1:W(1,0) TC2:W(1,0)

*CKT:CD 0 +D 0 0603C0.ckt FOOTPRINT

*FP:DRAW:xfig ATF3A.fig show
*calc:Layout 


SET:SAVEDATA true
.ends