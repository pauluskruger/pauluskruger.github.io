subck Opt2 0

R:Ri 0 1 r=50 temp=0 vac=2

SET:TEMP TEMP=290
SET:Q Q=50 $TEMP

CKT:I1 0 1 i1 i2 i3 I5C.ckt FOOTPRINT

CKT:S1 0 +i1 e1 S7C.ckt FOOTPRINT
CKT:S2 0 +i2 e2 S7C.ckt FOOTPRINT
CKT:U1 0 e1 e2 U1 i3 U5C.ckt FOOTPRINT

R:Ru 0 U1 r=50 temp=0
A:AD 0 U1 0 UD rin=1e6 rout=50 A=1e3 PW=1.2 PHASE=3.1416
SETPARAM:POWER-SCALE RI:R RU:R

FP:EQ:Q1 1 U1 ANG=0

SET:OPTI+I1: TI0:LEN(2.5e-3,5e-3) TI0:W(0.9e-3,2e-3) TI1:LEN(0.2e-3,5e-3) L0:L1:1(1,48) L1:L1:1(1,48) L2:L1:1(1,48,1) TG1:LEN(0.5e-3,2e-3) TG2:LEN(0.5e-3,2e-3) TI3:LEN(0.5e-3,5e-3) TI2:LEN(0.5e-3,5e-3) TI4:LEN(0.5e-3,5e-3) TFB:LEN(12e-3,20e-3) TFB2:LEN(2e-3,20e-3) TFB:W(0.3e-3,2e-3) TFB2:W(0.3e-3,2e-3) RFB:R1:R(1e1,1e5) TI1:W(0.5e-3,1e-3)  TG1:W(0.5e-3,1e-3) TG2:W(0.5e-3,1e-3)  TI2:W(0.5e-3,1e-3) TI3:W(0.7e-3,1e-3) TI4:W(0.7e-3,1e-3)
*  L3:L1:1(1,48,1)
*FUNC:F1 type=0 v1=1e-3 v2=1e-4 U1:TD1:LEN(1,1) U1:TD2:LEN(1,0)
SET:OPTU1 LD1:L1:1(1,48,1) LD2:L1:1(1,48,1) LU1:L1:1(1,48,1) LU2:L1:1(1,48,1) LU3:L1:1(1,48,1) LE1:L1:1(1,48,1) LE3:L1:1(1,48,1)
*SET:OPTU2 CD1:C1:1(1,10,1) CD2:C1:1(1,10,1) CUT:C1:1(1,41,1) CU:C1:1(1,41,1) CE1:C1:1(1,41,1) 
SET:OPTU2 CUT:C1:1(1,41,1) CU:C1:1(1,41,1) CE1:C1:1(1,41,1) 
SET:OPTU3 RUT:R1:R(1,100) RT2:R1:R(1,150) RFB:R1:R(1,1e3) RE1:R1:R(1,120) RE2:R1:R(1,1e5) RE3:R1:R(1,120)
*SET:OPTU4 TD1:LEN(0.5e-3,5e-3) TD2:LEN(0.5e-3,5e-3) TU1:LEN(0.5e-3,5e-3) TU2:LEN(0.5e-3,5e-3) TU3:LEN(0.5e-3,5e-3) TU4:LEN(0.5e-3,5e-3) 
SET:OPTU4 TU1:LEN(0.5e-3,2e-3) TU2:LEN(0.5e-3,5e-3) TU3:LEN(0.5e-3,5e-3) TU4:LEN(0.5e-3,5e-3)  F1:1(0.5e-3,2e-3) F1:2(0.1e-3,2.0e-3)
SET:OPTU5 TD1:W(0.3e-3,0.9e-3)   TD2:W(0.3e-3,0.9e-3)   TU1:W(0.3e-3,0.9e-3)   TU2:W(0.3e-3,0.9e-3)   TU3:W(0.3e-3,0.9e-3)   TU4:W(0.3e-3,0.9e-3)   
SET:OPTU+U1: $OPTU1 $OPTU2 $OPTU3 $OPTU4 $OPTU5 TU0:LEN(2.5e-3,5e-3) TU0:W(0.9e-3,2e-3)

set:OPT $OPTI $OPTU AD:PW(0.4,2)

LOADPARAM: Opt2U.dat $OPT
LOADPARAM: Opt3U.dat $OPT
LOADPARAM: O5C.dat $OPT



SET:OPTL1+I1:  FP:TFB:ANG(-90,90)   FP:TFB2:ANG(-40,40) FP:TG1:ANG(-50,30) FP:TG2:ANG(-30,30) FP:TI1:ANG(-30,30) FP:TI2:ANG(-30,30) FP:TI3:ANG(-30,30) FP:TI4:ANG(-30,30)
SET:OPTLS1+S1: FP:TD1:ANG(-60,-60) FP:TG2:ANG(-100,100) 
SET:OPTLS2+S2: FP:TD1:ANG(-100,100) FP:TG2:ANG(-100,100)
SET:OPTLU+U1: FP:TD2:ANG(-30,30) FP:TU1:ANG(0.1,0.1)  FP:TU2:ANG(-50,10)  FP:TU3:ANG(-50,10)  FP:TU3:ANG(-50,10) FP:TU4:ANG(-10,10) FP:TU0:ANG(-90,90)
SET:OPTL $OPTL1 $OPTLS1 $OPTLS2 $OPTLU
SET:FC1 F1=Layout:1 AVG1=1 WGH1=1e3
SET:FC2 F2=Layout:2 AVG2=1 WGH2=5
SET:FC3 F3=Layout:4 AVG3=1 WGH3=1

SET:FC $FC1 $FC2 $FC3

LOADPARAM: O5CL.dat $OPTL


set:OPSET dir=-1 START=1e9 STOP=1e9 STEP=0.1e9 maxsteps=10 savevar=O5CL.dat $FC $OPTL toll=1e-4

optim:step2 $OPSET
optim:rand $OPSET
optim:rands $OPSET P1=0.5 P2=2000
optim:step2 $OPSET
optim:rand $OPSET
optim:step2 $OPSET
optim:rand $OPSET
optim:step2 $OPSET
optim:rand $OPSET
optim:step2 $OPSET
optim:rand $OPSET
optim:step2 $OPSET
optim:rand $OPSET
optim:step2 $OPSET
optim:rand $OPSET

FP:DRAW:xfig O5CL.fig show
calc:Layout 
.ends
