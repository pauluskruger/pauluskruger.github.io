subck U2B 0 1 2 3 4
#include NN.subs

CKT:LD1 0 +1 h1 0603L0.ckt FOOTPRINT
CKT:LD2 0 +2 h2 0603L0.ckt FOOTPRINT

TMS:TD1 0 h1 a1c $DUR len=2e-3 w=0.3e-3 FOOTPRINT
TMS:TD2 0 h2 a2c $DUR len=2e-3 w=0.3e-3 ANG=-1 FOOTPRINT

TMS:TU1 0 a0 a1a $DUR len=2e-3 w=0.3e-3 ANG=-1 FOOTPRINT
TMS:TU2 0 a1b a1d $DUR len=2e-3 w=0.3e-3 ANG=-1 FOOTPRINT
TMS:TU3 0 a1e a2a $DUR len=2e-3 w=0.3e-3 ANG=-1 FOOTPRINT
TMS:TU4 0 a2b a3  $DUR len=2e-3 w=0.3e-3 ANG=-1  FOOTPRINT

*TMSTEE:TEE1 0 a1b a1a a1c M1=TU2 M2=TU1 M3=TD1 FOOTPRINT
TMSTEE:TEE1 0 a1c a1b a1a M1=TD1 M2=TU2 M3=TU1 FOOTPRINT
TMSTEE:TEE2 0 a2b a2a a2c M1=TU4 M2=TU3 M3=TD2 FOOTPRINT

CKT:RUT 0 -rt rt2 0603R0.ckt FOOTPRINT
CKT:RT2 0 rt3 rt2 rt4 0603RPS.ckt FOOTPRINT
CKT:CT2 0 rt4     0603CV.ckt FOOTPRINT
SETPARAM: CT2:C1:1 41
CKT:CUT 0 -rt3    0603CV.ckt FOOTPRINT

*CKT:LU1 0 +a0 rt 0603L0.ckt FOOTPRINT
CKT:LU1 0 -a0 ax rt 0603LPS.ckt FOOTPRINT
CKT:LU2 0 +a1d a1e 0603L0.ckt FOOTPRINT
CKT:LU3 0 +a3  P1 0603L0.ckt FOOTPRINT
CKT:CU  0 P1 P2  0603C0.ckt FOOTPRINT

CKT:RG1 0 P3 P2 R1 0603RPS.ckt FOOTPRINT
SETPARAM: RG1:R1:R 1e6 
TMSCNR:TCNR2 0 R1 +R1B $DUR w=0.9e-3 FOOTPRINT

CKT:RG2 0 +R1B R2 0603R0.ckt FOOTPRINT
SETPARAM: RG2:R1:R 1e6 
VIA:V2 0 R2 $DURVIA D=0.5e-3 FOOTPRINT


CKT:S3  0 +P3 U0 ATF3A.ckt FOOTPRINT
CKT:RFB 0 +U0 U1 U5 0603RPS.ckt FOOTPRINT

CKT:RE3 0 -U3b U9 0603R0.ckt FOOTPRINT
CKT:LE3 0 +U9 U10 0603L0.ckt FOOTPRINT
CKT:CE4 0 U10 0603CV.ckt FOOTPRINT
SETPARAM: CE4:C1:1 41

CKT:LE1 0 +U1 U2 0603L0.ckt FOOTPRINT
CKT:CE1 0 -U3c U4 0603C0.ckt FOOTPRINT
CKT:RE1 0 +U2 -U3 0603R0.ckt FOOTPRINT

TMSTEE:TEE3 0 -U3b +U3c +U3 M1=RE3:TP0 M2=CE1:TP0 M3=RE1:TP3   FOOTPRINT

CKT:RE2 0 U4 OUT 0603RVP.ckt FOOTPRINT

TMS:TU0 0 OUT 3 $DUR w=0.9e-3 len=2.5e-3 ANG=0.1 FOOTPRINT


CKT:CE2 0 U5 U6 0603C0.ckt FOOTPRINT
CKT:RE4 0 U6 4 0603RVP.ckt FOOTPRINT
SETPARAM: RE4:R1:R 1e6
SETPARAM: CE2:C1:1 41

FUNC:F1 type=0 v1=1e-3 v2=1e-4 TD1:LEN(1,1) TD2:LEN(1,0)

*FP:DRAW:xfig U5C.fig show
*calc:Layout 
.ends