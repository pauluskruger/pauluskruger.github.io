subck I2B 0 1 2 3 4 
#include NN.subs

TMS:TI0 0 1 in $DUR w=0.9e-3 len=2.5e-3 FOOTPRINT
CKT:L0 0 +in a5 0603L0.ckt FOOTPRINT
TMS:TI1 0 a5 a0a $DUR len=2e-3 w=0.9e-3 ANG=1 FOOTPRINT
*tee
TMS:TI2 0 a0b a0c $DUR len=1e-3 w=0.9e-3 ANG=1 FOOTPRINT
CKT:L1 0 +a0c a0d 0603L0.ckt FOOTPRINT
TMS:TI3 0 a0d a1a $DUR len=1e-3 w=0.9e-3 ANG=1 FOOTPRINT
*tee
TMS:TI4 0 a1b a1c $DUR len=1e-3 w=0.9e-3 ANG=1 FOOTPRINT
CKT:RFB 0 +a1c a7  0603R0.ckt FOOTPRINT
TMSCNR:TCNR1 0 a7 a2 $DUR w=0.9e-3 FOOTPRINT

TMS:TG1 0 b1 2 $DUR len=2e-3 w=0.9e-3 ANG=-10 FOOTPRINT
TMS:TG2 0 b2 3 $DUR len=2e-3 w=0.9e-3 ANG=-10 FOOTPRINT

TMSTEE:TEE1 0 a0b b1 a0a M1=TI2 M2=TG1 M3=TI1 FOOTPRINT
TMSTEE:TEE2 0 a1a a1b b2 M1=TI3 M2=TI4 M3=TG2 FOOTPRINT

TMS:TFB 0 a2 a3 $DUR len=1e-3 w=0.3e-3 ANG=20 FOOTPRINT

CKT:L2 0 +a3 fb 0603L0.ckt FOOTPRINT

TMS:TFB2 0 fb 4 $DUR len=14e-3 w=0.3e-3 ANG=20 FOOTPRINT

*FP:DRAW:xfig I5C.fig show
*calc:Layout 

.ends