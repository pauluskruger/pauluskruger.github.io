subck ATF35143CKT 0
#include NN.subs
SET:INVERT true
R:R1 0 A r=100 vac=2 temp=0
L:L1 A 1 l=10e-9 Q=50 temp=290  
CKT:S1     0 1 2 S7B.ckt FOOTPRINT
R:R2 0 2 r=200 temp=0

SETPARAM:POWER-SCALE R1:r R2:r

** Optimize function **
SET:FC1 F1=S1:M4:0:mag 		AVG1=1 		WGH1=1e0	START1=0.5e9	STOP1=1.8e9
SET:FC2 F2=S1:K        		AVG2=21	EX2=1.0	WGH2=1e4	START2=3e9
SET:FC3 F3=S1:Y:11:Re  		AVG3=21	EX3=1e-3	WGH3=1e6
SET:FC4 F4=S1:Y:22:Re  		AVG4=21	EX4=0	WGH4=1e5	START4=1e9
SET:FC5 F5=S1:K        		AVG5=21	EX5=1.2	WGH5=1e4	START5=5e9
SET:FC6 F6=S1:Y:11:Re		AVG6=21	EX6=0.02	WGH6=1e4	START6=0.5e9 STOP6=0.6e9

SET:FC $FC1 $FC2 $FC3 $FC4 $FC5 
*$FC6
** Optimize variables **
SET:OPT   S1:RD2:R1:R(1,100)  S1:TC2:LEN(1e-3,10e-3) S1:TC2:W(1e-3,2e-3) S1:TG2:LEN(1e-3,20e-3) S1:TG2:W(0.1e-3,2e-3) S1:TG1:LEN(1e-3,20e-3) S1:TG1:W(0.1e-3,2e-3) S1:TD1:LEN(0.1e-3,5e-3) S1:TD1:W(0.1e-3,2e-3) S1:CG1:C1:1(1,40,1) S1:RP1:R1:R(1,50) S1:LP1:L1:1(30,48,1) S1:T1:CGDV:1(1,10,1) S1:RP2:R1:R(1,200)
* S1:LG2:L(10e-9,50e-9) S1:R2:R1:R(1,50)

*  S1:S2:RD:R1:R(1,5000) 
*S1:C2:C(1e-13,1e-8)  
*S1:CS1V:1(1,41,1) S1:CS2V:1(1,41,1) S1:CS3V:1(1,41,1) S1:CS4V:1(1,41,1)
*SET:OPT S1:RD:R1:R(20,2000) S1:FL:1(0.1e-3,2e-3) S1:FW:1(0.05e-3,5e-3)
* S1:CD:C1:1(1,41)
*SET:OPT FL:1(0.11e-4,20e-3) FW:1(0.1e-3,5e-3) 
*RC:C1:1(1,30) * S1:TD:LEN(0.7e-3,3e-3)

LOADPARAM: S7Bo.dat  $OPT
SETPARAM: S1:T1:CGDV:1 1
*SETPARAM: S1:LP1:L1:1 48

** Optimize **
SET:OPSET dir=-1 start=0.1e9 stop=18.0011e9 step=0.1e9 maxsteps=0 savevar=S7Bo.dat $FC $OPT
optim:step2 $OPSET
*optim:rands $OPSET P1=0.8 P2=2000
*optim:step2 $OPSET
*optim:rand $OPSET
*optim:step2 $OPSET
*optim:rand $OPSET
*optim:step2 $OPSET

FP:DRAW:xfig S7Bo.fig show
calc:Layout 
*.ends

plot:"plots/S7B_K" freq S1:K
plot:"plots/S7B_Y" freq S1:Y:11:RE S1:Y:22:RE
calc:AC start=0.1e9 stop=18e9 step=0.1e9
CLOSEPRINT:

** plots **
SET:SIMFREQ start=0.05e9 stop=2.0e9 step=0.05e9

** Plots
plot:"plots/S7B_M.txt" freq S1:M4:0:mag S1:T1:M4:0:mag S1:T2:M4:0:mag 
*temp:2
*S1:S1:M4:0:mag S1:S1:T2:M4:0:mag
plot:"plots/S7B_N.txt" freq S1:AM4:0:db 
*gain:2:db
calc:AC $SIMFREQ
CLOSEPRINT:
.ends

