subck Sparm S G D

T:TA S G D atf35143i.s2p
.ends