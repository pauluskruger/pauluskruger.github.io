subck ATF35 0 1 2
#include NN.subs
SET:SAVEDATA true

CKT:T1 0 1 -D FET2.ckt FOOTPRINT

*CKT:CD 0 D D0 V1 0603CPS.ckt FOOTPRINT
*SETPARAM: CD:C1:1 1
*VIA:V1 0 V1 $DURVIA D=0.5e-3 FOOTPRINT

TMS:TD1 0 D X0 $DUR len=2e-3 w=0.3e-3 ANG=-50 FOOTPRINT


TMS:TC2 0 L L1 $DUR len=5e-3 w=1e-3 ang=-90 FOOTPRINT
*CKT:R2 0 L1 L2 0603R0.ckt FOOTPRINT
*TMS:TC3 0 L2 L3 $DUR len=5e-3 w=1e-3 FOOTPRINT

TMS:TG1 0 X1 X5 $DUR len=2e-3 w=0.4e-3 FOOTPRINT

TMSTEE:TEE1 0 X0 X1 L M1=TD1 M2=TG1 M3=TC2 FOOTPRINT

CKT:RP1 0 X2 X5 P1 0603RPS.ckt FOOTPRINT
CKT:LP1 0 +P1 -P2 0603L0.ckt FOOTPRINT

TMSCNR:TCNR1 0 +P2 -P2B $DUR w=0.9e-3 type=0 FOOTPRINT

CKT:RP2 0 +P2B P3 0603R0.ckt FOOTPRINT
CKT:CP1 0 P3 P4 0603C0.ckt FOOTPRINT
VIA:VP1 0 P4 $DURVIA D=0.5e-3 FOOTPRINT


CKT:CG1 0 X2 X3 0603C0.ckt FOOTPRINT

*DC on gate 2
CKT:RG1 0 X4 X3 -R1 0603RPS.ckt FOOTPRINT
SETPARAM: RG1:R1:R 1e6 
TMSCNR:TCNR2 0 +R1 -R1B   $DUR w=0.9e-3 FOOTPRINT

CKT:RG2 0 +R1B R2 0603R0.ckt FOOTPRINT
SETPARAM: RG2:R1:R 1e6 
VIA:V2 0 R2 $DURVIA D=0.5e-3 FOOTPRINT


TMS:TG2 0 X4 G2 $DUR len=1e-3 w=0.4e-3 ANG=-50 FOOTPRINT

CKT:T2 0 +G2 D2 ATF3A.ckt FOOTPRINT

CKT:RD2 0 D2 2 0603R0.ckt FOOTPRINT

SET:OPT  RD2:R1:R(1,500) TC2:LEN(1e-3,10e-3) TC2:W(1e-3,2e-3) TG2:LEN(1e-3,20e-3) TG2:W(0.1e-3,2e-3) TG1:LEN(1e-3,20e-3) TG1:W(0.1e-3,2e-3) TD1:LEN(0.1e-3,5e-3) TD1:W(0.1e-3,2e-3) CG1:C1:1(1,40,1) RP1:R1:R(1,50) LP1:L1:1(30,48,1) RP2:R1:R(1,200) T1:CGDV:1(1,10,1)
LOADPARAM: S7Bo2.dat  $OPT

*FP:DRAW:xfig S3.fig show
*calc:Layout 

.ends