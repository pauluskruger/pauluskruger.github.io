subck 0603C0 0 1 2 3 4

#include NN.subs

TMS:TP0 0 +1 +A1 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT
TMS:TP1 0 +2 -A1 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT

TMS:TP2 0 +4 +B1 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT
TMS:TP3 0 +3 -B1 $DUR len=0.45e-3 w=0.6e-3 FOOTPRINT

C:Cp A1 B1 c=0.01e-12

*TMSGAP:TG1 0 A2 B2 M1=TP1 M2=TP2



VIA:V1 0 B1 $DURVIA D=0.5e-3 FOOTPRINT="RPAD=0.01e-3"

TMSR:R1 0 A1 B1 $DURR W=0.9e-3 LEN=1.5e-3 R=100 $DISCRETE

FP:M2PADM:P A1 B1 D=0.9e-3 B=0.6e-3 W=0.9e-3 DIR1=1 DIR2=1 LABEL=R VALUE=R1:R

